OP AMP INTEGRATOR - SQUARE INPUT

.include LF356.MOD
XU1 3 2 7 4 6 LF356/NS

Vin 10 0 pulse(-1v 1v 0 0 0 1ms 2ms)

Rin 10 2 1kOhm
R1 3 0 0
Rf 2 6 1kohm
Cf 2 6 1uF
Vcc 7 0 9v
Vdd 4 0 -9v


.tran 1us 10ms
.control
run
plot v(10) v(6)
set xbrushwidth = 3
.endc
.end