HIGH PASS FILTER USING OP AMP

.include LF356.MOD
XU1 3 6 7 4 6 LF356/NS

Vin 10 0 dc=0 ac=1
c1 10 3 15.915nF
r1 3 0 10kOhm

vcc 7 0 15v
vee 4 0 -15v

.control
ac dec 100 1 1Meg
plot vdb(6)
set xbrushwidth=4
.endc
.end