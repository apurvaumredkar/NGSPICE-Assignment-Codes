OP AMP INTEGRATOR - SINE INPUT

.include LF356.MOD
XU1 3 2 7 4 6 LF356/NS

Vin 10 0 sine(0v 1v 1kHz)

Rin 10 2 1kOhm
R1 3 0 0
Rf 2 6 100kohm
Cf 2 6 1uF
Vcc 7 0 9v
Vdd 4 0 -9v


.tran 1us 10ms
.control
run
plot v(10) v(6)
set xbrushwidth = 3
.endc
.end

