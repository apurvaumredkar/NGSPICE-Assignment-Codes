BJT Amplifier
Vin 2 0 SINE(0V 0.01V 60Hz)
C1 1 2 10uF
Vcc 3 0 DC 5V
R1 1 3 68kOhm
Q1 5 1 0 mybjt
R2 1 0 10kOhm
R3 5 3 10kOhm
C2 5 6 10uF
Rload 6 0 100kOhm

.model mybjt npn(Is = 1e-15)
.tran 10us 50ms
.control
run
plot v(2) v(6)
set Xbrushwidth=4
.endc
.end