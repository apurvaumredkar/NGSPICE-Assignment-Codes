HALF ADDER USING CMOS

.model mosn nmos
.model mosp pmos

Va a 0 pulse(0 5 0 0 0 50ms 100ms)
Vb b 0 pulse(0 5 0 0 0 100ms 200ms)

.subckt xor a b z
vcc 1 0 dc 5v
m1 1 a s 1 mosp
m2 s a 0 0 mosn
m3 a b z 1 mosp
m4 z b s 0 mosn
.ends

.subckt and a b z
vcc 3 0 dc 5v
m1 4 a 3 3 mosp
m2 4 b 3 3 mosp
m3 5 a 4 0 mosn
m4 0 b 5 0 mosn
m5 z 4 3 3 mosp
m6 0 4 z 0 mosn
.ends

x3 a b sum xor
x4 a b carry and

.tran 100us 200ms
.control
run
plot v(a) v(b)+15 v(sum)+30 v(carry)+45
set xbrushwidth=4
.endc
.end
