NON INVERTING SUMMER

.include LF356.MOD
XU1 3 2 7 4 6 LF356/NS

V1 1 0 pulse(-2 2 0 0 0 50m 100m)
V2 10 0 pulse(-3 3 0 0 0 50m 100m)

R1 1 3 1k
R2 10 3 1k
Ra 2 0 1k
Rb 2 6 1k

vcc 7 0 15v
vee 4 0 -15v
.tran 10u 500m
.control
run
plot v(1) v(10) v(6)
.endc
.end