INVERTING SUMMER

.include LF356.MOD
XU1 0 2 7 4 6 LF356/NS

V1 1 0 pulse(-2 2 0 0 0 50ms 100ms)
V2 10 0 pulse(-3 3 0 0 0 50ms 100ms)

R1 1 2 1kOhm
R2 10 2 1kOhm
R3 2 6 1kOhm

vcc 7 0 15v
vee 4 0 -15v


.tran 10us 500ms
.control
run
plot v(1) v(10) v(6)
.endc
.end
