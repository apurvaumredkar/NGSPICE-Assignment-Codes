OSCILLATOR

R1 1 0 10kOhm
C1 1 2 1nF
R2 2 0 10kOhm
C2 2 3 1nF
R3 3 0 10kOhm
C3 3 5 1nF
R4 1 4 57kOhm
R5 5 4 6.8kOhm
Vcc 4 0 DC 10V
Q1 5 1 6 mybjt
R6 6 0 1.5kOhm
C4 6 0 0.1uF

.model mybjt npn(Is=1e-15)
.tran 10us 5ms
.control
run
plot v(4) v(5)
set Xbrushwidth=2
.endc
.end