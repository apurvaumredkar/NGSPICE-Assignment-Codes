BAND STOP FILTER USING OP AMP

.include LF356.MOD

XU1 3 6 7 4 6 LF356/NS
XU2 31 61 7 4 61 LF356/NS
XU3 32 22 7 4 62 LF356/NS

Vin 10 0 dc=0 ac=1

r1 10 3 10kOhm
c1 3 0 16nF

c2 10 31 1.6nF
r2 31 0 10kOhm


r3 6 22 10kOhm
r4 61 22 10kOhm
r5 22 62 10kOhm
r6 32 0 0 

vcc 7 0 15v
vee 4 0 -15v

.control
ac dec 100 1 1Meg
plot vdb(62) 
.endc
.end