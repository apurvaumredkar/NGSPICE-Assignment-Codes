Boolean Expression A+B+C
Va 1 0 PULSE(-5 5 0 0 0 50ns 100ns)
Vb 2 0 PULSE(-5 5 0 0 0 100ns 200ns)
Vc 3 0 PULSE(-5 5 0 0 0 200ns 400ns)

R1 4 2 10kOhm
Q1 5 4 6 mybjt
R2 7 3 10kOhm
Q2 5 7 6 mybjt
R3 6 0 10kOhm
Vcc 5 0 DC 5V

R4 8 6 10kOhm
Q3 5 8 9 mybjt
R5 10 1 10kOhm
Q4 5 10 9 mybjt
R6 9 0 10kOhm

.model mybjt npn(Is = 1e-15)
.tran 0.1NS 1000NS
.control
run
plot v(1) v(2)+15 v(3)+30 v(9)+45
.endc
.end