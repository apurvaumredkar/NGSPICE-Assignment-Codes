colpitt's oscillator

vcc 4 0 dc 12v

.model mybjt npn (is=1e-15)

q1 2 1 3 mybjt
r1 4 1 380kohm
rc 4 2 4.8kohm
cin 1 6 0.1uf
r2 1 0 72kohm
re 3 0 1.5kohm
ce 3 0 0.1uf

c1 2 0 10nf
c2 0 6 5nf
l1 2 6 100mh

.tran 0.01us 2.5ms

.control
run
plot v(4) v(2)
set xbrushwidth = 2
.endc
.end