NEGATIVE LEVEL TRIGGERED D FLIP FLOP

.model mosn nmos
.model mosp pmos

.subckt	nand	A	B	OP
Vdd 	1 	0 	dc 	5v 
m1 	1 	A 	OP 	1 	mosp
m2 	1 	B 	OP	1 	mosp 
m3 	OP 	A 	3 	0 	mosn
m4 	3 	B 	0 	0 	mosn
.ends

Vd	d	0	pulse(0 5 0 0 0 100ns 300ns)
Vclk	clk	0	pulse(0 5 0 0 0 125ns 250ns)

X1	d	d 	notd	nand
X2	d	clk	p1	nand
X3	notd	clk 	p2	nand
X4	p1	notq	q	nand
X5	p2	q	notq	nand

.tran 	1ns	1000ns
.control
run
plot	v(d)	v(clk)+10	v(q)+20	v(notq)+30
.endc
.end