BAND PASS FILTER USING OP AMP

.include LF356.MOD

XU1 3 6 7 4 6 LF356/NS
XU2 31 61 7 4 61 LF356/NS

Vin 10 0 dc=0 ac=1

c1 10 3 15.915nF
r1 3 0 10kOhm

r2 6 31 10kOhm
c2 31 0 0.053nF

vcc 7 0 15v
vee 4 0 -15v

.control
ac dec 10 1 10Meg
plot vdb(61)
.endc
.end